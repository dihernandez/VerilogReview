module hello_world();

	initial begin
		@$display("\n\t Hello World!\n");
	end
endmodule : hello_world